module decoder(
    input [31:0] instruction
);

endmodule